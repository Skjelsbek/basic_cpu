library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity stepper_motor_controller is
    Port
    (
        clk: in std_logic;
        dir: in std_logic; -- Direction
        JA: out std_logic_vector(3 downto 0); -- Outputs to coils on stepper motor
        dir_out: out std_logic
    );
end stepper_motor_controller;

architecture smc_arch of stepper_motor_controller is

    constant max_count: integer := 160000*2;
    constant control_level: integer := 79999*2+1;
    signal count: integer := 0;
    signal divided_clk: std_logic := '0';

    signal step: integer := 0;
    signal step_next: integer;
    signal test: std_logic;

begin

    counting: process (clk)
    begin
        if (rising_edge(clk)) then
            if (count < max_count) then
                count <= count + 1;
            else
                count <= 0;
            end if;
        end if;
    end process;

    pulsing: process (clk)
    begin
        if (rising_edge(clk)) then
            if (control_level > count) then
                divided_clk <= '0';
            else
                divided_clk <= '1';
            end if;
        end if;
    end process;

    update_state: process (divided_clk)
    begin
        if (rising_edge(divided_clk)) then
            step <= step_next;
        end if;
    end process;

    next_state_logic: process (step, dir)
    begin    
        case (step) is
            when 0 =>
                JA(0) <= '1';
                JA(1) <= '0';
                JA(2) <= '0';
                JA(3) <= '1';
            when 1 =>
                JA(0) <= '1';
                JA(1) <= '1';
                JA(2) <= '0';
                JA(3) <= '0';
            when 2 =>
                JA(0) <= '0';
                JA(1) <= '1';
                JA(2) <= '1';
                JA(3) <= '0';
            when 3 =>
                JA(0) <= '0';
                JA(1) <= '0';
                JA(2) <= '1';
                JA(3) <= '1';
            when others =>
                JA(0) <= '0';
                JA(1) <= '0';
                JA(2) <= '0';
                JA(3) <= '0';                                                                                                  
        end case;
            
        if (dir = '0') then
            if (step = 3) then
                step_next <= 0;
            else      
                step_next <= step + 1;                              
            end if;
        else
            if (step = 0) then
                step_next <= 3;                               
            else
                step_next <= step - 1;                            
            end if;
            
        end if;                 
    end process;
    dir_out <= dir;
end smc_arch;
